//-----------------------------------------------------------------------------
//
// Title       : TutorVHDL_tb_tim
// Design      : TutorVHDL
// Author      : KE
// Company     : AGH
//
//-----------------------------------------------------------------------------
//
// File        : TutorVHDL_TB_tim.v
// Generated   : Thu Nov 28 10:41:15 2019
// From        : C:\My_Designs\TutorVHDL_Cz0935\TutorVHDL\src\TestBench\TutorVHDL_TB_tim_settings.txt
// By          : tb_verilog.pl ver. ver 1.2s
//
//-----------------------------------------------------------------------------
//
// Description : 
//
//-----------------------------------------------------------------------------

`timescale 1ps / 1ps
module top_tb_tim;


//Internal signals declarations:

reg CLK;
reg CLR;
reg DataIn; 
wire DataOut;
reg LRCK_o;
reg MCLK;
reg SCLK_o; 
reg LOAD_o;
//reg LOW_ENABLE;
reg MID_ENABLE;
//reg HIGH_ENABLE;

// Unit Under Test port map
	Top UUT (
		.DataIn(DataIn),
		.DataOut(DataOut),
		.LRCK_o(LRCK_o),
		.CLR(CLR),
		.CLK(CLK),
		.MCLK(MCLK),
		.LOAD_o(LOAD_o),
		//.LOW_ENABLE(LOW_ENABLE),
		.MID_ENABLE(MID_ENABLE),
		//.HIGH_ENABLE(HIGH_ENABLE),
		.SCLK_o(SCLK_o));
		 
initial
	$monitor($realtime,,"ps %h %h %h %h %h %h %h %h %h",DataIn,DataOut,LRCK_o,CLR,CLK,MCLK,SCLK_o, LOAD_o, MID_ENABLE, );

//Below code was generated based on waveform file: "C:\My_Designs\TutorVHDL_Cz0935\TutorVHDL\compile\TutorVHDL.ver"

initial
begin : STIMUL // begin of stimulus process
	#0
	DataIn = 1'b1;
	CLR = 1'b1;
	CLK = 1'b0;	
    #5000; //0
	CLK = 1'b1;
    #5000; //50000
	CLR = 1'b0;
	CLK = 1'b0;
    #5000; //100000
	CLK = 1'b1;
    #5000; //150000
	CLR = 1'b1;
	CLK = 1'b0;
    #5000; //200000
	CLK = 1'b1;
    #5000; //250000
	CLK = 1'b0;
    #5000; //300000
	CLK = 1'b1;
    #5000; //350000
	CLK = 1'b0;
    #5000; //400000
	CLK = 1'b1;
    #5000; //450000
	CLK = 1'b0;
    #5000; //500000
	CLK = 1'b1;
    #5000; //550000
	CLK = 1'b0;
    #5000; //600000
	CLK = 1'b1;
    #5000; //650000
	CLK = 1'b0;
    #5000; //700000
	CLK = 1'b1;
    #5000; //750000
	CLK = 1'b0;
    #5000; //800000
	CLK = 1'b1;
    #5000; //850000
	CLK = 1'b0;
    #5000; //900000
	CLK = 1'b1;
    #5000; //950000   
	CLK = 1'b0;
    #5000; //1000000
	CLK = 1'b1;
    #5000; //1050000
	CLK = 1'b0;
    #25000; //1100000
	CLR = 1'b1;
    #25000; //1125000
	CLK = 1'b1;
    #5000; //1150000  
	CLK = 1'b0;
    #25000; //1200000
	CLR = 1'b0;
    #2500; //1225000
	CLK = 1'b1;
    #5000; //1250000
	CLK = 1'b0;
    #5000; //1300000
	CLK = 1'b1;
    #5000; //1350000
	CLK = 1'b0;		
    #5000; //1400000
	CLK = 1'b1;
    #5000; //1450000 
	CLK = 1'b0;		
    #5000; //1500000
	CLK = 1'b1;
    #5000; //1550000 
	CLK = 1'b0;
    #5000; //1600000
	CLK = 1'b1;
    #5000; //1650000
	CLK = 1'b0;
	#5000; //1700000
	CLK = 1'b1;
    #5000; //1750000 
	CLK = 1'b0;		
    #5000; //1800000
	CLK = 1'b1;
    #5000; //1850000
	CLK = 1'b0;
    #5000; //1900000
	CLK = 1'b1;
    #5000; //1950000
	CLK = 1'b0;
    #5000; //2000000
	CLK = 1'b1;	  
	DataIn = 1'b0;
    #5000; //2050000
	CLK = 1'b0;
    #5000; //2100000
	CLK = 1'b1;
    #5000; //2150000
	CLK = 1'b0;
    #5000; //2200000
	CLK = 1'b1;
    #5000; //2250000
	CLK = 1'b0;
    #5000; //2300000
	CLK = 1'b1;
    #5000; //2350000
	CLK = 1'b0;
    #5000; //2400000
	CLK = 1'b1;
    #5000; //2450000
	CLK = 1'b0;
    #5000; //2500000
	CLK = 1'b1;		 
	DataIn = 1'b1;
    #5000; //2550000
	CLK = 1'b0;
    #5000; //2600000
	CLK = 1'b1;
    #5000; //2650000
	CLK = 1'b0;
    #5000; //2700000
	CLK = 1'b1;		
	DataIn = 1'b0;
    #5000; //2750000
	CLK = 1'b0;
    #5000; //2800000
	CLK = 1'b1;
    #5000; //2850000
	CLK = 1'b0;
    #5000; //2900000
	CLK = 1'b1;
    #5000; //2950000
	CLK = 1'b0;
    #5000; //3000000
	CLK = 1'b1;
    #5000; //3050000
	CLK = 1'b0;
    #5000; //3100000
	CLK = 1'b1;
    #5000; //3150000
	CLK = 1'b0;
    #5000; //3200000
	CLK = 1'b1;
    #5000; //3250000
	CLK = 1'b0;
    #5000; //3300000
	CLK = 1'b1;
    #5000; //3350000
	CLK = 1'b0;
    #5000; //3400000
	CLK = 1'b1;
    #2500; //3450000
    #2500; //3475000
	CLK = 1'b0;
    #5000; //3500000
	CLK = 1'b1;		 
	DataIn = 1'b1;
    #5000; //3550000
	CLK = 1'b0;
    #5000; //3600000
	CLK = 1'b1;
    #5000; //3650000
	CLK = 1'b0;
    #5000; //3700000
	CLK = 1'b1;
    #5000; //3750000
	CLK = 1'b0;
    #5000; //3800000
	CLK = 1'b1;
    #5000; //3850000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;	
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
    #5000; //3900000
	CLK = 1'b1;
    #5000; //3950000
	CLK = 1'b0;
end // end of stimulus process
	



endmodule
